import top_pkg::*;

module top (
    input clk_sys_100MHz,
    input vga_hsync,
    input vga_vsync,
    input rgb444_t vga_rgb
  );
  
endmodule